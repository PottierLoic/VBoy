module main

const rom_types = [
	'ROM ONLY',
	'MBC1',
	'MBC1+RAM',
	'MBC1+RAM+BATTERY',
	'0x04 ???',
	'MBC2',
	'MBC2+BATTERY',
	'0x07 ???',
	'ROM+RAM 1',
	'ROM+RAM+BATTERY 1',
	'0x0A ???',
	'MMM01',
	'MMM01+RAM',
	'MMM01+RAM+BATTERY',
	'0x0E ???',
	'MBC3+TIMER+BATTERY',
	'MBC3+TIMER+RAM+BATTERY 2',
	'MBC3',
	'MBC3+RAM 2',
	'MBC3+RAM+BATTERY 2',
	'0x14 ???',
	'0x15 ???',
	'0x16 ???',
	'0x17 ???',
	'0x18 ???',
	'MBC5',
	'MBC5+RAM',
	'MBC5+RAM+BATTERY',
	'MBC5+RUMBLE',
	'MBC5+RUMBLE+RAM',
	'MBC5+RUMBLE+RAM+BATTERY',
	'0x1F ???',
	'MBC6',
	'0x21 ???',
	'MBC7+SENSOR+RUMBLE+RAM+BATTERY',
]

const lic_codes = [
	'None',
	'Nintendo R&D1',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Capcom',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Electronic Arts',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Hudson Soft',
	'b-ai',
	'kss',
	'Unknown',
	'pow',
	'Unknown',
	'PCM Complete',
	'san-x',
	'Unknown',
	'Unknown',
	'Kemco Japan',
	'seta',
	'Viacom',
	'Nintendo',
	'Bandai',
	'Ocean/Acclaim',
	'Konami',
	'Hector',
	'Unknown',
	'Taito',
	'Hudson',
	'Banpresto',
	'Unknown',
	'Ubi Soft',
	'Atlus',
	'Unknown',
	'Malibu',
	'Unknown',
	'angel',
	'Bullet-Proof',
	'Unknown',
	'irem',
	'Absolute',
	'Acclaim',
	'Activision',
	'American sammy',
	'Konami',
	'Hi tech entertainment',
	'LJN',
	'Matchbox',
	'Mattel',
	'Milton Bradley',
	'Titus',
	'Virgin',
	'Unknown',
	'Unknown',
	'LucasArts',
	'Unknown',
	'Unknown',
	'Ocean',
	'Unknown',
	'Electronic Arts',
	'Infogrames',
	'Interplay',
	'Broderbund',
	'sculptured',
	'Unknown',
	'sci',
	'Unknown',
	'Unknown',
	'THQ',
	'Accolade',
	'misawa',
	'Unknown',
	'Unknown',
	'lozc',
	'Unknown',
	'Unknown',
	'Tokuma Shoten Intermedia',
	'Tsukuda Original',
	'Unknown',
	'Unknown',
	'Unknown',
	'Chunsoft',
	'Video system',
	'Ocean/Acclaim',
	'Unknown',
	'Varie',
	"Yonezawa/s'pal",
	'Kaneko',
	'Unknown',
	'Pack in soft',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Unknown',
	'Konami (Yu-Gi-Oh!)',
]

const rom_sizes = [
	'32 KiB',
	'64 KiB',
	'128 KiB',
	'256 KiB',
	'512 KiB',
	'1 MiB',
	'2 MiB',
	'4 MiB',
	'8 MiB',
]

const ram_sizes = [
	'0',
	'-',
	'8 KiB',
	'32 KiB',
	'128 KiB',
	'64 KiB',
]
