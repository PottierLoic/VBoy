module main

import vboy

pub fn test_and() {

}