module vboy

pub fn (mut cpu Cpu) cpu_none() {
	println("test")
}
