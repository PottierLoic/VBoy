module vboy

type Cpu_fn_type = fn ()

fn (mut cpu Cpu) test_fn() {}

pub const cpu_fn = []

