module main

import vboy

fn main () {
	vboy.run()
}